/*
*  @file bsg_control_core.sv
*  @data March 2017
*  @brief Implementa a maquina de estados do BSG
**/

module bsg_control_core(


);







endmodule
