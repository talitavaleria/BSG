/*
*  @file modulator.svh
*  @data March 2017
*  @brief Implementa bsg TOP LEVEL
**/
module bsg(
);


  
endmodule
